`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:37:46 11/24/2017 
// Design Name: 
// Module Name:    Instruction_Memory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Instruction_Memory(
    input [31:0] a,
	 input CLK,
	 input WriteEnable,
	 input [5:0] keyboard,
    output reg [31:0] rd
    );
	 
	 reg [31:0] RAM[400:0];
	 
	 initial begin
	RAM[0] = 32'hE3A00002;
RAM[1] = 32'hE3A01000;
RAM[2] = 32'hE3A03000;
RAM[3] = 32'hE3A04000;
RAM[4] = 32'hE3A05004;
RAM[5] = 32'hE3A0A000;
RAM[6] = 32'hE3A0B0C0;
RAM[7] = 32'hE1A0B10B;
RAM[8] = 32'hE3A0C01A;
RAM[9] = 32'hE1A0C28C;
RAM[10] = 32'hE38CC01A;
RAM[11] = 32'hE1A0C38C;
RAM[12] = 32'hE58BC000;
RAM[13] = 32'hE3A0C000;
RAM[14] = 32'hEB0000d3;
RAM[15] = 32'hE2899000;
RAM[16] = 32'hE3A09000;
RAM[17] = 32'hE3590001;
RAM[18] = 32'h0Afffffb;
RAM[19] = 32'hE3A02001;
RAM[20] = 32'hEB000150;
RAM[21] = 32'hE352001E;
RAM[22] = 32'h1A0000b6;
RAM[23] = 32'hE1A08201;
RAM[24] = 32'hE2888002;
RAM[25] = 32'hE1A08108;
RAM[26] = 32'hE08AD008;
RAM[27] = 32'hE59D2000;
RAM[28] = 32'hE3520003;
RAM[29] = 32'h1A000016;
RAM[30] = 32'hE351000A;
RAM[31] = 32'h0B00006a;
RAM[32] = 32'hE35C0007;
RAM[33] = 32'h0A0000ed;
RAM[34] = 32'hE3A07004;
RAM[35] = 32'hEB0000cd;
RAM[36] = 32'hE3A02000;
RAM[37] = 32'hE1A02384;
RAM[38] = 32'hE1A08103;
RAM[39] = 32'hE08BD008;
RAM[40] = 32'hE59D4000;
RAM[41] = 32'hE2045070;
RAM[42] = 32'hE1A051A5;
RAM[43] = 32'hE1822005;
RAM[44] = 32'hE3844001;
RAM[45] = 32'hE58D4000;
RAM[46] = 32'hE28CC001;
RAM[47] = 32'hE1A0420C;
RAM[48] = 32'hE1822004;
RAM[49] = 32'hE1A0810C;
RAM[50] = 32'hE08BD008;
RAM[51] = 32'hE58D2000;
RAM[52] = 32'hEA0000c7;
RAM[53] = 32'hE3520005;
RAM[54] = 32'h1A000013;
RAM[55] = 32'hE351000A;
RAM[56] = 32'h0B000051;
RAM[57] = 32'hE35C0000;
RAM[58] = 32'h0A0000d4;
RAM[59] = 32'hE3A07004;
RAM[60] = 32'hEB0000b4;
RAM[61] = 32'hE3A02001;
RAM[62] = 32'hEB0000ef;
RAM[63] = 32'hEB0000fd;
RAM[64] = 32'hE08BD004;
RAM[65] = 32'hE59D5000;
RAM[66] = 32'hE2055001;
RAM[67] = 32'hE3550001;
RAM[68] = 32'h0A0000ca;
RAM[69] = 32'hEB000115;
RAM[70] = 32'hE3A02001;
RAM[71] = 32'hE3A07001;
RAM[72] = 32'hEB0000fe;
RAM[73] = 32'hE24CC001;
RAM[74] = 32'hEA0000b1;
RAM[75] = 32'hE352000D;
RAM[76] = 32'h1A000020;
RAM[77] = 32'hE351000A;
RAM[78] = 32'h0B00003b;
RAM[79] = 32'hE3A07004;
RAM[80] = 32'hEB0000a0;
RAM[81] = 32'hE3A02001;
RAM[82] = 32'hEB0000db;
RAM[83] = 32'hEB0000e9;
RAM[84] = 32'hE1A06005;
RAM[85] = 32'hE1A09004;
RAM[86] = 32'hE3A07007;
RAM[87] = 32'hEB000099;
RAM[88] = 32'hE3A02001;
RAM[89] = 32'hEB0000d4;
RAM[90] = 32'hE2052070;
RAM[91] = 32'hE1A021A2;
RAM[92] = 32'hE2067001;
RAM[93] = 32'hE1A06226;
RAM[94] = 32'hE1A06206;
RAM[95] = 32'hE1866007;
RAM[96] = 32'hE1866002;
RAM[97] = 32'hE3855001;
RAM[98] = 32'hE08BD009;
RAM[99] = 32'hE58D6000;
RAM[100] = 32'hE08BD008;
RAM[101] = 32'hE58D5000;
RAM[102] = 32'hE1A08103;
RAM[103] = 32'hE08BD008;
RAM[104] = 32'hE59D7000;
RAM[105] = 32'hE2079070;
RAM[106] = 32'hE3A02001;
RAM[107] = 32'hE3A07001;
RAM[108] = 32'hEB0000da;
RAM[109] = 32'hEA00008e;
RAM[110] = 32'hE3520004;
RAM[111] = 32'h1A000018;
RAM[112] = 32'hE351000A;
RAM[113] = 32'h0B000018;
RAM[114] = 32'hE1A08201;
RAM[115] = 32'hE2888004;
RAM[116] = 32'hE1A08108;
RAM[117] = 32'hE08AD008;
RAM[118] = 32'hE59D4000;
RAM[119] = 32'hE3540000;
RAM[120] = 32'h1A000008;
RAM[121] = 32'hE3530000;
RAM[122] = 32'h0A000094;
RAM[123] = 32'hE1A08003;
RAM[124] = 32'hE1A08108;
RAM[125] = 32'hE08BD008;
RAM[126] = 32'hE59D4000;
RAM[127] = 32'hE204400E;
RAM[128] = 32'hE1A030A4;
RAM[129] = 32'hEA00007a;
RAM[130] = 32'hE3A07004;
RAM[131] = 32'hEB00006d;
RAM[132] = 32'hE3A02000;
RAM[133] = 32'hEB0000a8;
RAM[134] = 32'hE2055070;
RAM[135] = 32'hE1A03225;
RAM[136] = 32'hEA000073;
RAM[137] = 32'hE352000C;
RAM[138] = 32'h1A000019;
RAM[139] = 32'hE3A04000;
RAM[140] = 32'hE1A08201;
RAM[141] = 32'hE0888004;
RAM[142] = 32'hE1A08108;
RAM[143] = 32'hE08AD008;
RAM[144] = 32'hE59D5000;
RAM[145] = 32'hE1A08104;
RAM[146] = 32'hE08AD008;
RAM[147] = 32'hE58D5000;
RAM[148] = 32'hE2844001;
RAM[149] = 32'hE3540010;
RAM[150] = 32'h1Afffff4;
RAM[151] = 32'hE3A04000;
RAM[152] = 32'hE3A05040;
RAM[153] = 32'hE3A06000;
RAM[154] = 32'hE08AD005;
RAM[155] = 32'hE58D6000;
RAM[156] = 32'hE2855004;
RAM[157] = 32'hE2844001;
RAM[158] = 32'hE35400B0;
RAM[159] = 32'h1Afffff9;
RAM[160] = 32'hE3A01001;
RAM[161] = 32'hE352000C;
RAM[162] = 32'h0A000046;
RAM[163] = 32'hE3A01000;
RAM[164] = 32'hE1A0F00E;
RAM[165] = 32'hE3520016;
RAM[166] = 32'h1A000023;
RAM[167] = 32'hE351000A;
RAM[168] = 32'h0Bffffe1;
RAM[169] = 32'hE2811001;
RAM[170] = 32'hE3A00000;
RAM[171] = 32'hE1A08103;
RAM[172] = 32'hE08BD008;
RAM[173] = 32'hE59D4000;
RAM[174] = 32'hE2044070;
RAM[175] = 32'hE1A04224;
RAM[176] = 32'hE3A05001;
RAM[177] = 32'hE1A08105;
RAM[178] = 32'hE08BD008;
RAM[179] = 32'hE59D6000;
RAM[180] = 32'hE206700E;
RAM[181] = 32'hE1A070A7;
RAM[182] = 32'hE1540007;
RAM[183] = 32'h1A00000e;
RAM[184] = 32'hE1A093A6;
RAM[185] = 32'hE1A062A9;
RAM[186] = 32'hE209901F;
RAM[187] = 32'hE1A08201;
RAM[188] = 32'hE0888000;
RAM[189] = 32'hE1A08108;
RAM[190] = 32'hE08AD008;
RAM[191] = 32'hE58D6000;
RAM[192] = 32'hE2800001;
RAM[193] = 32'hE1A08201;
RAM[194] = 32'hE0888000;
RAM[195] = 32'hE1A08108;
RAM[196] = 32'hE08AD008;
RAM[197] = 32'hE58D9000;
RAM[198] = 32'hE2800002;
RAM[199] = 32'hE2855001;
RAM[200] = 32'hE3550006;
RAM[201] = 32'h1Affffe6;
RAM[202] = 32'hEA00001e;
RAM[203] = 32'hE351000A;
RAM[204] = 32'h0Bffffbd;
RAM[205] = 32'hEA000041;
RAM[206] = 32'hE352001F;
RAM[207] = 32'h1A000009;
RAM[208] = 32'hE3500002;
RAM[209] = 32'h0Affff3c;
RAM[210] = 32'hE2400001;
RAM[211] = 32'hE1A08201;
RAM[212] = 32'hE0888000;
RAM[213] = 32'hE1A08108;
RAM[214] = 32'hE08AD008;
RAM[215] = 32'hE3A02000;
RAM[216] = 32'hE58D2000;
RAM[217] = 32'hEAffff34;
RAM[218] = 32'hE3500010;
RAM[219] = 32'h0Affff32;
RAM[220] = 32'hE1A08201;
RAM[221] = 32'hE0888000;
RAM[222] = 32'hE1A08108;
RAM[223] = 32'hE08AD008;
RAM[224] = 32'hE58D2000;
RAM[225] = 32'hE2800001;
RAM[226] = 32'hEAffff2b;
RAM[227] = 32'hE3A0201C;
RAM[228] = 32'hE08AD004;
RAM[229] = 32'hE58D2000;
RAM[230] = 32'hE3A0201D;
RAM[231] = 32'hE08AD005;
RAM[232] = 32'hE58D2000;
RAM[233] = 32'hE1A0F00E;
RAM[234] = 32'hE2811001;
RAM[235] = 32'hE3A00002;
RAM[236] = 32'hE1A08201;
RAM[237] = 32'hE1A08108;
RAM[238] = 32'hE1A04008;
RAM[239] = 32'hE2845004;
RAM[240] = 32'hEBfffff1;
RAM[241] = 32'hEAffff1c;
RAM[242] = 32'hE1A08201;
RAM[243] = 32'hE0888007;
RAM[244] = 32'hE1A08108;
RAM[245] = 32'hE08AD008;
RAM[246] = 32'hE59D4000;
RAM[247] = 32'hE1A04284;
RAM[248] = 32'hE2888004;
RAM[249] = 32'hE08AD008;
RAM[250] = 32'hE59D5000;
RAM[251] = 32'hE1844005;
RAM[252] = 32'hE1A0F00E;
RAM[253] = 32'hE2811001;
RAM[254] = 32'hE1A08201;
RAM[255] = 32'hE1A08108;
RAM[256] = 32'hE3A05004;
RAM[257] = 32'hE08AD008;
RAM[258] = 32'hE58D5000;
RAM[259] = 32'hE2888004;
RAM[260] = 32'hE3A0500F;
RAM[261] = 32'hE08AD008;
RAM[262] = 32'hE58D5000;
RAM[263] = 32'hE2888004;
RAM[264] = 32'hE3A0500E;
RAM[265] = 32'hE08AD008;
RAM[266] = 32'hE58D5000;
RAM[267] = 32'hE2888004;
RAM[268] = 32'hE3A05005;
RAM[269] = 32'hE08AD008;
RAM[270] = 32'hE58D5000;
RAM[271] = 32'hEAffffd9;
RAM[272] = 32'hE2811001;
RAM[273] = 32'hE1A08201;
RAM[274] = 32'hE1A08108;
RAM[275] = 32'hE3A05009;
RAM[276] = 32'hE08AD008;
RAM[277] = 32'hE58D5000;
RAM[278] = 32'hE2888004;
RAM[279] = 32'hE3A0500E;
RAM[280] = 32'hE08AD008;
RAM[281] = 32'hE58D5000;
RAM[282] = 32'hE2888004;
RAM[283] = 32'hE3A05016;
RAM[284] = 32'hE08AD008;
RAM[285] = 32'hE58D5000;
RAM[286] = 32'hE2888004;
RAM[287] = 32'hE3A05001;
RAM[288] = 32'hE08AD008;
RAM[289] = 32'hE58D5000;
RAM[290] = 32'hE2888004;
RAM[291] = 32'hE3A0500C;
RAM[292] = 32'hE08AD008;
RAM[293] = 32'hE58D5000;
RAM[294] = 32'hE2888004;
RAM[295] = 32'hE3A05009;
RAM[296] = 32'hE08AD008;
RAM[297] = 32'hE58D5000;
RAM[298] = 32'hE2888004;
RAM[299] = 32'hE3A05004;
RAM[300] = 32'hE08AD008;
RAM[301] = 32'hE58D5000;
RAM[302] = 32'hEAffffba;
RAM[303] = 32'hE1A08002;
RAM[304] = 32'hE1A08108;
RAM[305] = 32'hE08BD008;
RAM[306] = 32'hE59D5000;
RAM[307] = 32'hE1A073A5;
RAM[308] = 32'hE1570004;
RAM[309] = 32'hE3A07001;
RAM[310] = 32'h0A000003;
RAM[311] = 32'hE2822001;
RAM[312] = 32'hE3520008;
RAM[313] = 32'h1Afffff4;
RAM[314] = 32'hE3A07000;
RAM[315] = 32'hE3570000;
RAM[316] = 32'h0Affffd2;
RAM[317] = 32'hE1A0F00E;
RAM[318] = 32'hE1A04008;
RAM[319] = 32'hE1A08103;
RAM[320] = 32'hE08BD008;
RAM[321] = 32'hE59D7000;
RAM[322] = 32'hE2079070;
RAM[323] = 32'hE205700E;
RAM[324] = 32'hE1A07187;
RAM[325] = 32'hE1570009;
RAM[326] = 32'h1Affffc8;
RAM[327] = 32'hE1A0F00E;
RAM[328] = 32'hE1A08102;
RAM[329] = 32'hE08BD008;
RAM[330] = 32'hE59D6000;
RAM[331] = 32'hE206800E;
RAM[332] = 32'hE1A08188;
RAM[333] = 32'hE1580009;
RAM[334] = 32'h0A000003;
RAM[335] = 32'hE2822001;
RAM[336] = 32'hE3520008;
RAM[337] = 32'h1Afffff5;
RAM[338] = 32'hE3A07000;
RAM[339] = 32'hE3570000;
RAM[340] = 32'hE1A08103;
RAM[341] = 32'hE08BD008;
RAM[342] = 32'hE59D6000;
RAM[343] = 32'h1A000001;
RAM[344] = 32'hE1A060A6;
RAM[345] = 32'hE1A06086;
RAM[346] = 32'hE58D6000;
RAM[347] = 32'hE1A0F00E;
RAM[348] = 32'hE2847004;
RAM[349] = 32'hE08BD007;
RAM[350] = 32'hE59D6000;
RAM[351] = 32'hE08BD004;
RAM[352] = 32'hE58D6000;
RAM[353] = 32'hE2844004;
RAM[354] = 32'hE2822001;
RAM[355] = 32'hE3520008;
RAM[356] = 32'h1Afffff6;
RAM[357] = 32'hE1A0F00E;
RAM[358] = 32'hE3A04000;
RAM[359] = 32'hE3A05000;
RAM[360] = 32'hE3A06000;
RAM[361] = 32'hE3A07000;
RAM[362] = 32'hE3A08000;
RAM[363] = 32'hE3A09000;
RAM[364] = 32'hE288D000;
RAM[365] = 32'hE1A0F00E;
	end

	 always @(a)
		begin
			rd = RAM[a/4];
		end
	
	 always @(posedge CLK)
		begin
			if(WriteEnable)
				begin
					RAM[17] <= {{31'b1110001101011001000000000000000},keyboard[0]};
					RAM[19] <= {{27'b111000111010000000100000000},keyboard[5:1]};
				end
		end
	 
endmodule
