`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:37:46 11/24/2017 
// Design Name: 
// Module Name:    Instruction_Memory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Instruction_Memory(
    input [31:0] a,
	 input CLK,
	 input WriteEnable,
	 input [5:0] keyboard,
    output reg [31:0] rd
    );
	 
	 reg [31:0] RAM[400:0];
	 
	 initial begin

RAM[0] = 32'hE3A00002;
RAM[1] = 32'hE3A01000;
RAM[2] = 32'hE3A03000;
RAM[3] = 32'hE3A04000;
RAM[4] = 32'hE3A05004;
RAM[5] = 32'hE3A0AC00;
RAM[6] = 32'hE3A0BCC0;
RAM[7] = 32'hE3A0C000;
RAM[8] = 32'hEB0000f2;
RAM[9] = 32'hE3A09000;
RAM[10] = 32'hE3590001;
RAM[11] = 32'h1A000007;
RAM[12] = 32'hE3A02000;
RAM[13] = 32'hE1A07000;
RAM[14] = 32'hE1A08201;
RAM[15] = 32'hE0888007;
RAM[16] = 32'hE1A08108;
RAM[17] = 32'hE08AD008;
RAM[18] = 32'hE58D2000;
RAM[19] = 32'hEAfffff4;
RAM[20] = 32'hE3A0201E;
RAM[21] = 32'hE352001E;
RAM[22] = 32'h1A0000ce;
RAM[23] = 32'hE3A07002;
RAM[24] = 32'hE1A08201;
RAM[25] = 32'hE0888007;
RAM[26] = 32'hE1A08108;
RAM[27] = 32'hE08AD008;
RAM[28] = 32'hE59D2000;
RAM[29] = 32'hE3520003;
RAM[30] = 32'h1A000019;
RAM[31] = 32'hE351000A;
RAM[32] = 32'h0B000079;
RAM[33] = 32'hE35C0007;
RAM[34] = 32'h0A000109;
RAM[35] = 32'hE3A07004;
RAM[36] = 32'hEB0000e7;
RAM[37] = 32'hE3A02000;
RAM[38] = 32'hE1A02384;
RAM[39] = 32'hE1A08003;
RAM[40] = 32'hE1A08108;
RAM[41] = 32'hE08BD008;
RAM[42] = 32'hE59D4000;
RAM[43] = 32'hE2045070;
RAM[44] = 32'hE1A051A5;
RAM[45] = 32'hE1822005;
RAM[46] = 32'hE3844001;
RAM[47] = 32'hE08BD006;
RAM[48] = 32'hE58D4000;
RAM[49] = 32'hE28CC001;
RAM[50] = 32'hE1A0420C;
RAM[51] = 32'hE1822004;
RAM[52] = 32'hE1A0800C;
RAM[53] = 32'hE1A08108;
RAM[54] = 32'hE08BD008;
RAM[55] = 32'hE58D2000;
RAM[56] = 32'hEA0000de;
RAM[57] = 32'hE3520005;
RAM[58] = 32'h1A000020;
RAM[59] = 32'hE351000A;
RAM[60] = 32'h0B00005d;
RAM[61] = 32'hE35C0000;
RAM[62] = 32'h0A0000ed;
RAM[63] = 32'hE3A07004;
RAM[64] = 32'hEB0000cb;
RAM[65] = 32'hE3A02001;
RAM[66] = 32'hEB00010a;
RAM[67] = 32'hEB00011a;
RAM[68] = 32'hE08BD004;
RAM[69] = 32'hE59D5000;
RAM[70] = 32'hE2055070;
RAM[71] = 32'hEB000138;
RAM[72] = 32'hE3A02001;
RAM[73] = 32'hE3A07001;
RAM[74] = 32'hEB00011e;
RAM[75] = 32'hE3A09001;
RAM[76] = 32'hE1A08009;
RAM[77] = 32'hE1A08108;
RAM[78] = 32'hE08BD008;
RAM[79] = 32'hE59D7000;
RAM[80] = 32'hE207700E;
RAM[81] = 32'hE1A07187;
RAM[82] = 32'hE1570005;
RAM[83] = 32'hE1A04008;
RAM[84] = 32'hE1A02009;
RAM[85] = 32'h02499001;
RAM[86] = 32'h0A000129;
RAM[87] = 32'hE2899001;
RAM[88] = 32'hE3590007;
RAM[89] = 32'h1Afffff1;
RAM[90] = 32'hE24CC001;
RAM[91] = 32'hEA0000bb;
RAM[92] = 32'hE352000D;
RAM[93] = 32'h1A000022;
RAM[94] = 32'hE351000A;
RAM[95] = 32'h0B00003a;
RAM[96] = 32'hE3530000;
RAM[97] = 32'h0A0000ca;
RAM[98] = 32'hE3A07004;
RAM[99] = 32'hEB0000a8;
RAM[100] = 32'hE3A02000;
RAM[101] = 32'hEB0000e7;
RAM[102] = 32'hEB0000f7;
RAM[103] = 32'hE1A06005;
RAM[104] = 32'hE1A09004;
RAM[105] = 32'hE3A07008;
RAM[106] = 32'hEB0000a1;
RAM[107] = 32'hE3A02000;
RAM[108] = 32'hEB0000e0;
RAM[109] = 32'hE2052070;
RAM[110] = 32'hE206700F;
RAM[111] = 32'hE1A063A6;
RAM[112] = 32'hE1A06386;
RAM[113] = 32'hE1866007;
RAM[114] = 32'hE1866002;
RAM[115] = 32'hE3855001;
RAM[116] = 32'hE08BD009;
RAM[117] = 32'hE58D6000;
RAM[118] = 32'hE08BD008;
RAM[119] = 32'hE58D5000;
RAM[120] = 32'hE1A08003;
RAM[121] = 32'hE1A08108;
RAM[122] = 32'hE08BD008;
RAM[123] = 32'hE59D7000;
RAM[124] = 32'hE2079070;
RAM[125] = 32'hE3A02001;
RAM[126] = 32'hE3A07001;
RAM[127] = 32'hEB0000e9;
RAM[128] = 32'hEA000096;
RAM[129] = 32'hE3520004;
RAM[130] = 32'h1A000017;
RAM[131] = 32'hE351000A;
RAM[132] = 32'h0B000015;
RAM[133] = 32'hE3A07008;
RAM[134] = 32'hE1A08201;
RAM[135] = 32'hE0888007;
RAM[136] = 32'hE1A08108;
RAM[137] = 32'hE08AD008;
RAM[138] = 32'hE59D4000;
RAM[139] = 32'hE354001D;
RAM[140] = 32'h1A000006;
RAM[141] = 32'hE1A08003;
RAM[142] = 32'hE1A08108;
RAM[143] = 32'hE08AD008;
RAM[144] = 32'hE59D4000;
RAM[145] = 32'hE204400E;
RAM[146] = 32'hE1A030A4;
RAM[147] = 32'hEA000083;
RAM[148] = 32'hE3A07008;
RAM[149] = 32'hEB000076;
RAM[150] = 32'hE3A02001;
RAM[151] = 32'hEB0000b5;
RAM[152] = 32'hE2055070;
RAM[153] = 32'hE1A03225;
RAM[154] = 32'hEA00007c;
RAM[155] = 32'hE352000C;
RAM[156] = 32'h1A00001b;
RAM[157] = 32'hE3A02000;
RAM[158] = 32'hE1A07004;
RAM[159] = 32'hE1A08201;
RAM[160] = 32'hE0888007;
RAM[161] = 32'hE1A08108;
RAM[162] = 32'hE08AD008;
RAM[163] = 32'hE59D5000;
RAM[164] = 32'hE1A08004;
RAM[165] = 32'hE1A08108;
RAM[166] = 32'hE08AD008;
RAM[167] = 32'hE58D5000;
RAM[168] = 32'hE2844001;
RAM[169] = 32'hE3540010;
RAM[170] = 32'h1Afffff2;
RAM[171] = 32'hE3A04000;
RAM[172] = 32'hE3A05040;
RAM[173] = 32'hE3A06000;
RAM[174] = 32'hE08AD005;
RAM[175] = 32'hE58D6000;
RAM[176] = 32'hE2855004;
RAM[177] = 32'hE2844001;
RAM[178] = 32'hE35400B0;
RAM[179] = 32'h1Afffff9;
RAM[180] = 32'hE3A01001;
RAM[181] = 32'hE352000C;
RAM[182] = 32'h0A00004b;
RAM[183] = 32'hE3A01000;
RAM[184] = 32'hE1A0F00E;
RAM[185] = 32'hE3520016;
RAM[186] = 32'h1A000027;
RAM[187] = 32'hE351000A;
RAM[188] = 32'h0Bffffdd;
RAM[189] = 32'hE2811001;
RAM[190] = 32'hE3A00000;
RAM[191] = 32'hE1A08003;
RAM[192] = 32'hE1A08108;
RAM[193] = 32'hE08BD008;
RAM[194] = 32'hE59D4000;
RAM[195] = 32'hE2044070;
RAM[196] = 32'hE1A04224;
RAM[197] = 32'hE3A05001;
RAM[198] = 32'hE1A08005;
RAM[199] = 32'hE1A08108;
RAM[200] = 32'hE08BD008;
RAM[201] = 32'hE59D6000;
RAM[202] = 32'hE206700E;
RAM[203] = 32'hE1A070A7;
RAM[204] = 32'hE1540007;
RAM[205] = 32'h1A000010;
RAM[206] = 32'hE1A093A6;
RAM[207] = 32'hE1A062A9;
RAM[208] = 32'hE209900F;
RAM[209] = 32'hE1A07000;
RAM[210] = 32'hE1A08201;
RAM[211] = 32'hE0888007;
RAM[212] = 32'hE1A08108;
RAM[213] = 32'hE08AD008;
RAM[214] = 32'hE58D6000;
RAM[215] = 32'hE2800001;
RAM[216] = 32'hE1A07000;
RAM[217] = 32'hE1A08201;
RAM[218] = 32'hE0888007;
RAM[219] = 32'hE1A08108;
RAM[220] = 32'hE08AD008;
RAM[221] = 32'hE58D9000;
RAM[222] = 32'hE2800002;
RAM[223] = 32'hE2855001;
RAM[224] = 32'hE3550007;
RAM[225] = 32'h1Affffe3;
RAM[226] = 32'hEA00001f;
RAM[227] = 32'hE351000A;
RAM[228] = 32'h0Bffffb5;
RAM[229] = 32'hEA000046;
RAM[230] = 32'hE352001F;
RAM[231] = 32'h1A000009;
RAM[232] = 32'hE3500002;
RAM[233] = 32'h0Affff1e;
RAM[234] = 32'hE2400001;
RAM[235] = 32'hE1A07000;
RAM[236] = 32'hE1A08201;
RAM[237] = 32'hE0888007;
RAM[238] = 32'hE1A08108;
RAM[239] = 32'hE08AD008;
RAM[240] = 32'hE58D2000;
RAM[241] = 32'hEAffff16;
RAM[242] = 32'hE350000F;
RAM[243] = 32'h0Affff14;
RAM[244] = 32'hE1A07000;
RAM[245] = 32'hE1A08201;
RAM[246] = 32'hE0888007;
RAM[247] = 32'hE1A08108;
RAM[248] = 32'hE08BD008;
RAM[249] = 32'hE58D2000;
RAM[250] = 32'hE2800001;
RAM[251] = 32'hEAffff0c;
RAM[252] = 32'hE3A0201C;
RAM[253] = 32'hE08AD004;
RAM[254] = 32'hE58D2000;
RAM[255] = 32'hE3A0201D;
RAM[256] = 32'hE08AD005;
RAM[257] = 32'hE58D2000;
RAM[258] = 32'hE1A0F00E;
RAM[259] = 32'hE2811001;
RAM[260] = 32'hE3A00002;
RAM[261] = 32'hE3A07000;
RAM[262] = 32'hE1A08201;
RAM[263] = 32'hE0888007;
RAM[264] = 32'hE1A08108;
RAM[265] = 32'hE1A04008;
RAM[266] = 32'hE2845004;
RAM[267] = 32'hEBffffef;
RAM[268] = 32'hEAfffefb;
RAM[269] = 32'hE1A08201;
RAM[270] = 32'hE0888007;
RAM[271] = 32'hE1A08108;
RAM[272] = 32'hE08AD008;
RAM[273] = 32'hE59D4000;
RAM[274] = 32'hE1A04284;
RAM[275] = 32'hE2888004;
RAM[276] = 32'hE08AD008;
RAM[277] = 32'hE59D5000;
RAM[278] = 32'hE1844005;
RAM[279] = 32'hE1A0F00E;
RAM[280] = 32'hE2811001;
RAM[281] = 32'hE3A07000;
RAM[282] = 32'hE1A08201;
RAM[283] = 32'hE0888007;
RAM[284] = 32'hE1A08108;
RAM[285] = 32'hE3A05004;
RAM[286] = 32'hE08AD008;
RAM[287] = 32'hE58D5000;
RAM[288] = 32'hE2888004;
RAM[289] = 32'hE3A0500F;
RAM[290] = 32'hE08AD008;
RAM[291] = 32'hE58D5000;
RAM[292] = 32'hE2888004;
RAM[293] = 32'hE3A0500E;
RAM[294] = 32'hE08AD008;
RAM[295] = 32'hE58D5000;
RAM[296] = 32'hE2888004;
RAM[297] = 32'hE3A05005;
RAM[298] = 32'hE08AD008;
RAM[299] = 32'hE58D5000;
RAM[300] = 32'hEAffffd5;
RAM[301] = 32'hE2811001;
RAM[302] = 32'hE3A07000;
RAM[303] = 32'hE1A08201;
RAM[304] = 32'hE0888007;
RAM[305] = 32'hE1A08108;
RAM[306] = 32'hE3A05009;
RAM[307] = 32'hE08AD008;
RAM[308] = 32'hE58D5000;
RAM[309] = 32'hE2888004;
RAM[310] = 32'hE3A0500E;
RAM[311] = 32'hE08AD008;
RAM[312] = 32'hE58D5000;
RAM[313] = 32'hE2888004;
RAM[314] = 32'hE3A05016;
RAM[315] = 32'hE08AD008;
RAM[316] = 32'hE58D5000;
RAM[317] = 32'hE58D5000;
RAM[318] = 32'hE2888004;
RAM[319] = 32'hE3A05001;
RAM[320] = 32'hE08AD008;
RAM[321] = 32'hE58D5000;
RAM[322] = 32'hE2888004;
RAM[323] = 32'hE3A0500C;
RAM[324] = 32'hE08AD008;
RAM[325] = 32'hE58D5000;
RAM[326] = 32'hE2888004;
RAM[327] = 32'hE3A05009;
RAM[328] = 32'hE08AD008;
RAM[329] = 32'hE58D5000;
RAM[330] = 32'hE2888004;
RAM[331] = 32'hE3A05004;
RAM[332] = 32'hE08AD008;
RAM[333] = 32'hE58D5000;
RAM[334] = 32'hEAffffb4;
RAM[335] = 32'hE1A08002;
RAM[336] = 32'hE1A08108;
RAM[337] = 32'hE08BD008;
RAM[338] = 32'hE59D5000;
RAM[339] = 32'hE1A073A5;
RAM[340] = 32'hE1A07387;
RAM[341] = 32'hE1A04384;
RAM[342] = 32'hE1570004;
RAM[343] = 32'hE3A07001;
RAM[344] = 32'h0A000003;
RAM[345] = 32'hE2822001;
RAM[346] = 32'hE15C0002;
RAM[347] = 32'h1Afffff2;
RAM[348] = 32'hE3A07000;
RAM[349] = 32'hE3570000;
RAM[350] = 32'h0Affffce;
RAM[351] = 32'hE1A0F00E;
RAM[352] = 32'hE1A04008;
RAM[353] = 32'hE1A08003;
RAM[354] = 32'hE1A08108;
RAM[355] = 32'hE08BD008;
RAM[356] = 32'hE59D7000;
RAM[357] = 32'hE2079070;
RAM[358] = 32'hE205700E;
RAM[359] = 32'hE1A07187;
RAM[360] = 32'hE1570009;
RAM[361] = 32'h1Affffc3;
RAM[362] = 32'hE1A0F00E;
RAM[363] = 32'hE1A08002;
RAM[364] = 32'hE1A08108;
RAM[365] = 32'hE08BD008;
RAM[366] = 32'hE59D6000;
RAM[367] = 32'hE206800E;
RAM[368] = 32'hE1A08188;
RAM[369] = 32'hE1580009;
RAM[370] = 32'h0A000003;
RAM[371] = 32'hE2822001;
RAM[372] = 32'hE3520007;
RAM[373] = 32'h1Afffff4;
RAM[374] = 32'hE3A07000;
RAM[375] = 32'hE3570000;
RAM[376] = 32'hE1A08003;
RAM[377] = 32'hE1A08108;
RAM[378] = 32'hE08BD008;
RAM[379] = 32'hE59D6000;
RAM[380] = 32'h1A000001;
RAM[381] = 32'hE1A060A6;
RAM[382] = 32'hE1A06086;
RAM[383] = 32'hE08BD008;
RAM[384] = 32'hE58D6000;
RAM[385] = 32'hE1A0F00E;
RAM[386] = 32'hE2847004;
RAM[387] = 32'hE08BD007;
RAM[388] = 32'hE59D6000;
RAM[389] = 32'hE08BD004;
RAM[390] = 32'hE58D6000;
RAM[391] = 32'hE2844004;
RAM[392] = 32'hE2822001;
RAM[393] = 32'hE3520007;
RAM[394] = 32'h1Afffff6;
RAM[395] = 32'hE1A0F00E;
	end

	 always @(a)
		begin
			rd = RAM[a/4];
		end
	
	 always @(negedge CLK)
		begin
			if(WriteEnable)
				begin
					RAM[9] <= {{31'b1110001101011001000000000000000},keyboard[0]};
					RAM[6] <= {{27'b111000111010000000100000000},keyboard[5:1]};
				end
		end
	 
endmodule
