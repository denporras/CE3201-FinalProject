`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:22:44 11/20/2017 
// Design Name: 
// Module Name:    TopLevelModule 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module TopLevelModule(
    );

	wire [3:0] A1;
   wire [3:0] A2;
   wire [3:0] A3;
   wire [31:0] WD3;
	wire [31:0] R15;
	wire	WE3;
   wire [31:0] RD1;
   wire [31:0] RD2;
	wire CLK;

	


endmodule
